module webcam_desktop

import openpnp_capture

#flag -I @VMODROOT/c
